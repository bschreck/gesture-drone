library verilog;
use verilog.vl_types.all;
entity Gest_Rec_test is
end Gest_Rec_test;
