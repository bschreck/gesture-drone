library verilog;
use verilog.vl_types.all;
entity Hover_test is
end Hover_test;
