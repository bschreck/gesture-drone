`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:13:29 12/01/2014 
// Design Name: 
// Module Name:    Display 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Display(
    input clock,
    input reset,
    input [15:0] x1,
    input [15:0] y1,
	 input [15:0] z1,
	 input [15:0] x2,
	 input [15:0] y2,
	 input [15:0] z2
    );


endmodule
