library verilog;
use verilog.vl_types.all;
entity On_FSM_test is
end On_FSM_test;
